module Ctrl(
	input [5:0] opcode;
	output RegDst, Branch, MemtoReg, MemWrite, ALUSrc, RegWrite;
	output [1:0] ALUOp;
);

module  Registers(
    input [5:0] read_reg1, read_reg2, write_reg;
    input reg_write;
    input [31:0] write_data;
    output [31:0] read_data1, read_data2;
);

assign read_data1 = read_data2 = 32'd0;

endmodule
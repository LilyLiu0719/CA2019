module ALU32(
	
);
